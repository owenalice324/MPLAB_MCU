library verilog;
use verilog.vl_types.all;
entity cpu_test is
end cpu_test;
